module uart_fifo_buffer(CLOCK_TX, CLOCK_RX, RESET, SEND, LOAD_FIFO, READ_FIFO, READ_BUFF, DATA_IN_FIFO,
		NINTO, NINTI, LD_FIFO_DONE, RD_FIFO_DONE, DATA_OUT_BUFF);
input CLOCK_TX, CLOCK_RX, RESET, SEND, LOAD_FIFO, READ_FIFO, READ_BUFF;
input [7:0] DATA_IN_FIFO;
output NINTO, NINTI, LD_FIFO_DONE, RD_FIFO_DONE;
output [7:0] DATA_OUT_BUFF;

wire [7:0] DATA_OUT_FIFO, DATA_OUT_UART;

fifo inst_fifo_tx(CLOCK_TX, RESET, LOAD_FIFO, READ_FIFO, DATA_IN_FIFO, LD_FIFO_DONE, RD_FIFO_DONE, DATA_OUT_FIFO);
uart inst_uart(CLOCK_TX, CLOCK_RX, RESET, SEND, DATA_OUT_FIFO, NINTO, NINTI, DATA_OUT_UART);
buffer_rx inst_buffer_rx(CLOCK_RX, RESET, READ_BUFF, DATA_OUT_UART, DATA_OUT_BUFF);

endmodule